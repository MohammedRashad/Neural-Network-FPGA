library IEEE; 
use IEEE.STD_LOGIC_1164.all; 

package package_types is 

type INT_ARRAY is array (integer range <>) of integer;
type matrix is array (integer range <>, integer range <>) of integer;

end package_types; 


package body package_types is 


end package_types; 
